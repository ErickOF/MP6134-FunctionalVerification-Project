// Based on: https://www.edaplayground.com/x/Yk4N
class scoreboard;
  logic [31:0] instruction_queue [$];
  logic [31:0] data_queue [$];
endclass : scoreboard
