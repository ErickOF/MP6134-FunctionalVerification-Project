typedef enum logic [6:0] {
  r_type = 7'b011_0011;
  i_type = 7'b001_0011; //TODO: only for: ADDI, XORI, ORI, ANDI, SLLI, SRLI, SRAI, SLTI and SLTIU
  s_type = 7'b010_0011;
  b_type = 7'b110_0011;
  u_type = 7'b001_0111; //TODO: only for AUIPC
  j_type = 7'b110_1111; //TODO: only for JAL
} inst_type_e;