// Based on: https://www.edaplayground.com/x/Yk4N
interface dut_intf(input clk);
endinterface : dut_intf
