// Based on: https://www.edaplayground.com/x/Yk4N
class stimulus;
endclass : stimulus
