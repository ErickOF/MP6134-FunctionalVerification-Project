`ifndef _RISCV_ITEMS_PKG_SV_
`define _RISCV_ITEMS_PKG_SV_

package riscv_items_pkg;

  import uvm_pkg::*;

  `include "riscv_input_item.svh"
  `include "riscv_output_item.svh"

endpackage : riscv_items_pkg

`endif // _RISCV_ITEMS_PKG_SV_