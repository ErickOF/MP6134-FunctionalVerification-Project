interface darksimv_hdl_xtor(input CLK);

  

endinterface : darksimv_hdl_xtor
