// Based on: https://www.edaplayground.com/x/Yk4N
class scoreboard;
endclass : scoreboard
